entity readout_complete_simple_top is
  port (
    
  ) ;
end entity;


architecture arch of readout_complete_simple_top is

    

begin

    

end architecture ;